library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM is
port (CLK : in std_logic;
      EN : in std_logic;
      ADDR : in std_logic_vector(9 downto 0);
      DATA : out std_logic_vector(7 downto 0));
end ROM;

architecture syn of ROM is
    type rom_type is array (1023 downto 0) of std_logic_vector (7 downto 0);                 
    signal ROM : rom_type:= (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00");
    
	 signal rdata : std_logic_vector(7 downto 0);
begin

    rdata <= ROM(conv_integer(ADDR));

    process (CLK)
    begin
        if (CLK'event and CLK = '1') then
            if (EN = '1') then
                DATA <= rdata;
				else
					DATA <= "ZZZZZZZZ";
            end if;
        end if;
    end process;

end syn;

				