----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:52:41 06/05/2016 
-- Design Name: 
-- Module Name:    mem_control - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mem_control is
	port(
				IR: in std_logic_vector(7 downto 0);
				CONT: in std_logic_vector(2 downto 0);
				salida_mem_control : out std_logic_vector(24 downto 0)
			);
end mem_control;

architecture Behavioral of mem_control is

	signal se�ales_de_control : std_logic_vector(27 downto 0);

begin

	se�ales_de_control <= X"0050100" WHEN IR&CONT = "00000000000" ELSE
          X"0004000" WHEN IR&CONT = "00000000001" ELSE
          X"0802000" WHEN IR&CONT = "00000000010" ELSE
          X"0050100" WHEN IR&CONT = "00000001000" ELSE
          X"0004000" WHEN IR&CONT = "00000001001" ELSE
          X"0802001" WHEN IR&CONT = "00000001010" ELSE
          X"0050100" WHEN IR&CONT = "00000010000" ELSE
          X"0004000" WHEN IR&CONT = "00000010001" ELSE
          X"0802002" WHEN IR&CONT = "00000010010" ELSE
          X"0050100" WHEN IR&CONT = "00000011000" ELSE
          X"0004000" WHEN IR&CONT = "00000011001" ELSE
          X"0050100" WHEN IR&CONT = "00000011010" ELSE
          X"0008000" WHEN IR&CONT = "00000011011" ELSE
          X"0802003" WHEN IR&CONT = "00000011100" ELSE
          X"0050100" WHEN IR&CONT = "00000100000" ELSE
          X"0004000" WHEN IR&CONT = "00000100001" ELSE
          X"0801004" WHEN IR&CONT = "00000100010" ELSE
          X"0050100" WHEN IR&CONT = "00000101000" ELSE
          X"0004000" WHEN IR&CONT = "00000101001" ELSE
          X"0801005" WHEN IR&CONT = "00000101010" ELSE
          X"0050100" WHEN IR&CONT = "00000110000" ELSE
          X"0004000" WHEN IR&CONT = "00000110001" ELSE
          X"0801006" WHEN IR&CONT = "00000110010" ELSE
          X"0050100" WHEN IR&CONT = "00000111000" ELSE
          X"0004000" WHEN IR&CONT = "00000111001" ELSE
          X"0050100" WHEN IR&CONT = "00000111010" ELSE
          X"0008000" WHEN IR&CONT = "00000111011" ELSE
          X"0801007" WHEN IR&CONT = "00000111100" ELSE
          X"0050100" WHEN IR&CONT = "00001000000" ELSE
          X"0004000" WHEN IR&CONT = "00001000001" ELSE
          X"0800808" WHEN IR&CONT = "00001000010" ELSE
          X"0050100" WHEN IR&CONT = "00001001000" ELSE
          X"0004000" WHEN IR&CONT = "00001001001" ELSE
          X"0800809" WHEN IR&CONT = "00001001010" ELSE
          X"0050100" WHEN IR&CONT = "00001010000" ELSE
          X"0004000" WHEN IR&CONT = "00001010001" ELSE
          X"080080A" WHEN IR&CONT = "00001010010" ELSE
          X"0050100" WHEN IR&CONT = "00001011000" ELSE
          X"0004000" WHEN IR&CONT = "00001011001" ELSE
          X"0050100" WHEN IR&CONT = "00001011010" ELSE
          X"0008000" WHEN IR&CONT = "00001011011" ELSE
          X"080080B" WHEN IR&CONT = "00001011100" ELSE
          X"0050100" WHEN IR&CONT = "00010011000" ELSE
          X"0004000" WHEN IR&CONT = "00010011001" ELSE
          X"0050100" WHEN IR&CONT = "00010011010" ELSE
          X"0008000" WHEN IR&CONT = "00010011011" ELSE
          X"0010020" WHEN IR&CONT = "00010011100" ELSE
          X"0008000" WHEN IR&CONT = "00010011101" ELSE
          X"0802003" WHEN IR&CONT = "00010011110" ELSE
          X"0050100" WHEN IR&CONT = "00011100000" ELSE
          X"0004000" WHEN IR&CONT = "00011100001" ELSE
          X"0050100" WHEN IR&CONT = "00011100010" ELSE
          X"0008000" WHEN IR&CONT = "00011100011" ELSE
          X"0010020" WHEN IR&CONT = "00011100100" ELSE
          X"0008010" WHEN IR&CONT = "00011100101" ELSE
          X"0800200" WHEN IR&CONT = "00011100110" ELSE
          X"0050100" WHEN IR&CONT = "00010111000" ELSE
          X"0004000" WHEN IR&CONT = "00010111001" ELSE
          X"0050100" WHEN IR&CONT = "00010111010" ELSE
          X"0008000" WHEN IR&CONT = "00010111011" ELSE
          X"0010020" WHEN IR&CONT = "00010111100" ELSE
          X"0008000" WHEN IR&CONT = "00010111101" ELSE
          X"0801007" WHEN IR&CONT = "00010111110" ELSE
          X"0050100" WHEN IR&CONT = "00011101000" ELSE
          X"0004000" WHEN IR&CONT = "00011101001" ELSE
          X"0050100" WHEN IR&CONT = "00011101010" ELSE
          X"0008000" WHEN IR&CONT = "00011101011" ELSE
          X"0010020" WHEN IR&CONT = "00011101100" ELSE
          X"0008015" WHEN IR&CONT = "00011101101" ELSE
          X"0800200" WHEN IR&CONT = "00011101110" ELSE
          X"0050100" WHEN IR&CONT = "00011011000" ELSE
          X"0004000" WHEN IR&CONT = "00011011001" ELSE
          X"0050100" WHEN IR&CONT = "00011011010" ELSE
          X"0008000" WHEN IR&CONT = "00011011011" ELSE
          X"0010020" WHEN IR&CONT = "00011011100" ELSE
          X"0008000" WHEN IR&CONT = "00011011101" ELSE
          X"080080B" WHEN IR&CONT = "00011011110" ELSE
          X"0050100" WHEN IR&CONT = "00011110000" ELSE
          X"0004000" WHEN IR&CONT = "00011110001" ELSE
          X"0050100" WHEN IR&CONT = "00011110010" ELSE
          X"0008000" WHEN IR&CONT = "00011110011" ELSE
          X"0010020" WHEN IR&CONT = "00011110100" ELSE
          X"000801A" WHEN IR&CONT = "00011110101" ELSE
          X"0800200" WHEN IR&CONT = "00011110110" ELSE
          X"0050100" WHEN IR&CONT = "0010----000" ELSE
          X"0004000" WHEN IR&CONT = "0010----001" ELSE
          X"0820000" WHEN IR&CONT = "0010----010" ELSE
          X"0050100" WHEN IR&CONT = "00110000000" ELSE
          X"0004000" WHEN IR&CONT = "00110000001" ELSE
          X"0882000" WHEN IR&CONT = "00110000010" ELSE
          X"0050100" WHEN IR&CONT = "00110001000" ELSE
          X"0004000" WHEN IR&CONT = "00110001001" ELSE
          X"0882001" WHEN IR&CONT = "00110001010" ELSE
          X"0050100" WHEN IR&CONT = "00110010000" ELSE
          X"0004000" WHEN IR&CONT = "00110010001" ELSE
          X"0882002" WHEN IR&CONT = "00110010010" ELSE
          X"0050100" WHEN IR&CONT = "00110011000" ELSE
          X"0004000" WHEN IR&CONT = "00110011001" ELSE
          X"0050100" WHEN IR&CONT = "00110011010" ELSE
          X"0008000" WHEN IR&CONT = "00110011011" ELSE
          X"0882003" WHEN IR&CONT = "00110011100" ELSE
          X"0050100" WHEN IR&CONT = "00110100000" ELSE
          X"0004000" WHEN IR&CONT = "00110100001" ELSE
          X"0881004" WHEN IR&CONT = "00110100010" ELSE
          X"0050100" WHEN IR&CONT = "00110101000" ELSE
          X"0004000" WHEN IR&CONT = "00110101001" ELSE
          X"0881005" WHEN IR&CONT = "00110101010" ELSE
          X"0050100" WHEN IR&CONT = "00110110000" ELSE
          X"0004000" WHEN IR&CONT = "00110110001" ELSE
          X"0881006" WHEN IR&CONT = "00110110010" ELSE
          X"0050100" WHEN IR&CONT = "00110111000" ELSE
          X"0004000" WHEN IR&CONT = "00110111001" ELSE
          X"0050100" WHEN IR&CONT = "00110111010" ELSE
          X"0008000" WHEN IR&CONT = "00110111011" ELSE
          X"0881007" WHEN IR&CONT = "00110111100" ELSE
          X"0050100" WHEN IR&CONT = "00111000000" ELSE
          X"0004000" WHEN IR&CONT = "00111000001" ELSE
          X"0880808" WHEN IR&CONT = "00111000010" ELSE
          X"0050100" WHEN IR&CONT = "00111001000" ELSE
          X"0004000" WHEN IR&CONT = "00111001001" ELSE
          X"0880809" WHEN IR&CONT = "00111001010" ELSE
          X"0050100" WHEN IR&CONT = "00111010000" ELSE
          X"0004000" WHEN IR&CONT = "00111010001" ELSE
          X"088080A" WHEN IR&CONT = "00111010010" ELSE
          X"0050100" WHEN IR&CONT = "00111011000" ELSE
          X"0004000" WHEN IR&CONT = "00111011001" ELSE
          X"0050100" WHEN IR&CONT = "00111011010" ELSE
          X"0008000" WHEN IR&CONT = "00111011011" ELSE
          X"088080B" WHEN IR&CONT = "00111011100" ELSE
          X"0050100" WHEN IR&CONT = "01000000000" ELSE
          X"0004000" WHEN IR&CONT = "01000000001" ELSE
          X"0902000" WHEN IR&CONT = "01000000010" ELSE
          X"0050100" WHEN IR&CONT = "01000001000" ELSE
          X"0004000" WHEN IR&CONT = "01000001001" ELSE
          X"0902001" WHEN IR&CONT = "01000001010" ELSE
          X"0050100" WHEN IR&CONT = "01000010000" ELSE
          X"0004000" WHEN IR&CONT = "01000010001" ELSE
          X"0902002" WHEN IR&CONT = "01000010010" ELSE
          X"0050100" WHEN IR&CONT = "01000011000" ELSE
          X"0004000" WHEN IR&CONT = "01000011001" ELSE
          X"0050100" WHEN IR&CONT = "01000011010" ELSE
          X"0008000" WHEN IR&CONT = "01000011011" ELSE
          X"0902003" WHEN IR&CONT = "01000011100" ELSE
          X"0050100" WHEN IR&CONT = "01000100000" ELSE
          X"0004000" WHEN IR&CONT = "01000100001" ELSE
          X"0901004" WHEN IR&CONT = "01000100010" ELSE
          X"0050100" WHEN IR&CONT = "01000101000" ELSE
          X"0004000" WHEN IR&CONT = "01000101001" ELSE
          X"0901005" WHEN IR&CONT = "01000101010" ELSE
          X"0050100" WHEN IR&CONT = "01000110000" ELSE
          X"0004000" WHEN IR&CONT = "01000110001" ELSE
          X"0901006" WHEN IR&CONT = "01000110010" ELSE
          X"0050100" WHEN IR&CONT = "01000111000" ELSE
          X"0004000" WHEN IR&CONT = "01000111001" ELSE
          X"0050100" WHEN IR&CONT = "01000111010" ELSE
          X"0008000" WHEN IR&CONT = "01000111011" ELSE
          X"0901007" WHEN IR&CONT = "01000111100" ELSE
          X"0050100" WHEN IR&CONT = "01001000000" ELSE
          X"0004000" WHEN IR&CONT = "01001000001" ELSE
          X"0900808" WHEN IR&CONT = "01001000010" ELSE
          X"0050100" WHEN IR&CONT = "01001001000" ELSE
          X"0004000" WHEN IR&CONT = "01001001001" ELSE
          X"0900809" WHEN IR&CONT = "01001001010" ELSE
          X"0050100" WHEN IR&CONT = "01001010000" ELSE
          X"0004000" WHEN IR&CONT = "01001010001" ELSE
          X"090080A" WHEN IR&CONT = "01001010010" ELSE
          X"0050100" WHEN IR&CONT = "01001011000" ELSE
          X"0004000" WHEN IR&CONT = "01001011001" ELSE
          X"0050100" WHEN IR&CONT = "01001011010" ELSE
          X"0008000" WHEN IR&CONT = "01001011011" ELSE
          X"090080B" WHEN IR&CONT = "01001011100" ELSE
          X"0050100" WHEN IR&CONT = "01010000000" ELSE
          X"0004000" WHEN IR&CONT = "01010000001" ELSE
          X"0902000" WHEN IR&CONT = "01010000010" ELSE
          X"0050100" WHEN IR&CONT = "01010001000" ELSE
          X"0004000" WHEN IR&CONT = "01010001001" ELSE
          X"0902001" WHEN IR&CONT = "01010001010" ELSE
          X"0050100" WHEN IR&CONT = "01010010000" ELSE
          X"0004000" WHEN IR&CONT = "01010010001" ELSE
          X"0902002" WHEN IR&CONT = "01010010010" ELSE
          X"0050100" WHEN IR&CONT = "01010011000" ELSE
          X"0004000" WHEN IR&CONT = "01010011001" ELSE
          X"0050100" WHEN IR&CONT = "01010011010" ELSE
          X"0008000" WHEN IR&CONT = "01010011011" ELSE
          X"0902003" WHEN IR&CONT = "01010011100" ELSE
          X"0050100" WHEN IR&CONT = "01010100000" ELSE
          X"0004000" WHEN IR&CONT = "01010100001" ELSE
          X"0901004" WHEN IR&CONT = "01010100010" ELSE
          X"0050100" WHEN IR&CONT = "01010101000" ELSE
          X"0004000" WHEN IR&CONT = "01010101001" ELSE
          X"0901005" WHEN IR&CONT = "01010101010" ELSE
          X"0050100" WHEN IR&CONT = "01010110000" ELSE
          X"0004000" WHEN IR&CONT = "01010110001" ELSE
          X"0901006" WHEN IR&CONT = "01010110010" ELSE
          X"0050100" WHEN IR&CONT = "01010111000" ELSE
          X"0004000" WHEN IR&CONT = "01010111001" ELSE
          X"0050100" WHEN IR&CONT = "01010111010" ELSE
          X"0008000" WHEN IR&CONT = "01010111011" ELSE
          X"0901007" WHEN IR&CONT = "01010111100" ELSE
          X"0050100" WHEN IR&CONT = "01011000000" ELSE
          X"0004000" WHEN IR&CONT = "01011000001" ELSE
          X"0900808" WHEN IR&CONT = "01011000010" ELSE
          X"0050100" WHEN IR&CONT = "01011001000" ELSE
          X"0004000" WHEN IR&CONT = "01011001001" ELSE
          X"0900809" WHEN IR&CONT = "01011001010" ELSE
          X"0050100" WHEN IR&CONT = "01011010000" ELSE
          X"0004000" WHEN IR&CONT = "01011010001" ELSE
          X"090080A" WHEN IR&CONT = "01011010010" ELSE
          X"0050100" WHEN IR&CONT = "01011011000" ELSE
          X"0004000" WHEN IR&CONT = "01011011001" ELSE
          X"0050100" WHEN IR&CONT = "01011011010" ELSE
          X"0008000" WHEN IR&CONT = "01011011011" ELSE
          X"090080B" WHEN IR&CONT = "01011011100" ELSE
          X"0050100" WHEN IR&CONT = "01100000000" ELSE
          X"0004000" WHEN IR&CONT = "01100000001" ELSE
          X"0A02000" WHEN IR&CONT = "01100000010" ELSE
          X"0050100" WHEN IR&CONT = "01100001000" ELSE
          X"0004000" WHEN IR&CONT = "01100001001" ELSE
          X"0A02001" WHEN IR&CONT = "01100001010" ELSE
          X"0050100" WHEN IR&CONT = "01100010000" ELSE
          X"0004000" WHEN IR&CONT = "01100010001" ELSE
          X"0A02002" WHEN IR&CONT = "01100010010" ELSE
          X"0050100" WHEN IR&CONT = "01100011000" ELSE
          X"0004000" WHEN IR&CONT = "01100011001" ELSE
          X"0050100" WHEN IR&CONT = "01100011010" ELSE
          X"0008000" WHEN IR&CONT = "01100011011" ELSE
          X"0A02003" WHEN IR&CONT = "01100011100" ELSE
          X"0050100" WHEN IR&CONT = "01100100000" ELSE
          X"0004000" WHEN IR&CONT = "01100100001" ELSE
          X"0A01004" WHEN IR&CONT = "01100100010" ELSE
          X"0050100" WHEN IR&CONT = "01100101000" ELSE
          X"0004000" WHEN IR&CONT = "01100101001" ELSE
          X"0A01005" WHEN IR&CONT = "01100101010" ELSE
          X"0050100" WHEN IR&CONT = "01100110000" ELSE
          X"0004000" WHEN IR&CONT = "01100110001" ELSE
          X"0A01006" WHEN IR&CONT = "01100110010" ELSE
          X"0050100" WHEN IR&CONT = "01100111000" ELSE
          X"0004000" WHEN IR&CONT = "01100111001" ELSE
          X"0050100" WHEN IR&CONT = "01100111010" ELSE
          X"0008000" WHEN IR&CONT = "01100111011" ELSE
          X"0A01007" WHEN IR&CONT = "01100111100" ELSE
          X"0050100" WHEN IR&CONT = "01101000000" ELSE
          X"0004000" WHEN IR&CONT = "01101000001" ELSE
          X"0A00808" WHEN IR&CONT = "01101000010" ELSE
          X"0050100" WHEN IR&CONT = "01101001000" ELSE
          X"0004000" WHEN IR&CONT = "01101001001" ELSE
          X"0A00809" WHEN IR&CONT = "01101001010" ELSE
          X"0050100" WHEN IR&CONT = "01101010000" ELSE
          X"0004000" WHEN IR&CONT = "01101010001" ELSE
          X"0A0080A" WHEN IR&CONT = "01101010010" ELSE
          X"0050100" WHEN IR&CONT = "01101011000" ELSE
          X"0004000" WHEN IR&CONT = "01101011001" ELSE
          X"0050100" WHEN IR&CONT = "01101011010" ELSE
          X"0008000" WHEN IR&CONT = "01101011011" ELSE
          X"0A0080B" WHEN IR&CONT = "01101011100" ELSE
          X"0050100" WHEN IR&CONT = "01110000000" ELSE
          X"0004000" WHEN IR&CONT = "01110000001" ELSE
          X"0A82000" WHEN IR&CONT = "01110000010" ELSE
          X"0050100" WHEN IR&CONT = "01110001000" ELSE
          X"0004000" WHEN IR&CONT = "01110001001" ELSE
          X"0A82001" WHEN IR&CONT = "01110001010" ELSE
          X"0050100" WHEN IR&CONT = "01110010000" ELSE
          X"0004000" WHEN IR&CONT = "01110010001" ELSE
          X"0A82002" WHEN IR&CONT = "01110010010" ELSE
          X"0050100" WHEN IR&CONT = "01110011000" ELSE
          X"0004000" WHEN IR&CONT = "01110011001" ELSE
          X"0050100" WHEN IR&CONT = "01110011010" ELSE
          X"0008000" WHEN IR&CONT = "01110011011" ELSE
          X"0A82003" WHEN IR&CONT = "01110011100" ELSE
          X"0050100" WHEN IR&CONT = "01110100000" ELSE
          X"0004000" WHEN IR&CONT = "01110100001" ELSE
          X"0A81004" WHEN IR&CONT = "01110100010" ELSE
          X"0050100" WHEN IR&CONT = "01110101000" ELSE
          X"0004000" WHEN IR&CONT = "01110101001" ELSE
          X"0A81005" WHEN IR&CONT = "01110101010" ELSE
          X"0050100" WHEN IR&CONT = "01110110000" ELSE
          X"0004000" WHEN IR&CONT = "01110110001" ELSE
          X"0A81006" WHEN IR&CONT = "01110110010" ELSE
          X"0050100" WHEN IR&CONT = "01110111000" ELSE
          X"0004000" WHEN IR&CONT = "01110111001" ELSE
          X"0050100" WHEN IR&CONT = "01110111010" ELSE
          X"0008000" WHEN IR&CONT = "01110111011" ELSE
          X"0A81007" WHEN IR&CONT = "01110111100" ELSE
          X"0050100" WHEN IR&CONT = "01111000000" ELSE
          X"0004000" WHEN IR&CONT = "01111000001" ELSE
          X"0A80808" WHEN IR&CONT = "01111000010" ELSE
          X"0050100" WHEN IR&CONT = "01111001000" ELSE
          X"0004000" WHEN IR&CONT = "01111001001" ELSE
          X"0A80809" WHEN IR&CONT = "01111001010" ELSE
          X"0050100" WHEN IR&CONT = "01111010000" ELSE
          X"0004000" WHEN IR&CONT = "01111010001" ELSE
          X"0A8080A" WHEN IR&CONT = "01111010010" ELSE
          X"0050100" WHEN IR&CONT = "01111011000" ELSE
          X"0004000" WHEN IR&CONT = "01111011001" ELSE
          X"0050100" WHEN IR&CONT = "01111011010" ELSE
          X"0008000" WHEN IR&CONT = "01111011011" ELSE
          X"0A8080B" WHEN IR&CONT = "01111011100" ELSE
          X"0050100" WHEN IR&CONT = "10000000000" ELSE
          X"0004000" WHEN IR&CONT = "10000000001" ELSE
          X"0B02040" WHEN IR&CONT = "10000000010" ELSE
          X"0050100" WHEN IR&CONT = "10000001000" ELSE
          X"0004000" WHEN IR&CONT = "10000001001" ELSE
          X"0B02041" WHEN IR&CONT = "10000001010" ELSE
          X"0050100" WHEN IR&CONT = "10000010000" ELSE
          X"0004000" WHEN IR&CONT = "10000010001" ELSE
          X"0B02042" WHEN IR&CONT = "10000010010" ELSE
          X"0050100" WHEN IR&CONT = "10000011000" ELSE
          X"0004000" WHEN IR&CONT = "10000011001" ELSE
          X"0050100" WHEN IR&CONT = "10000011010" ELSE
          X"0008000" WHEN IR&CONT = "10000011011" ELSE
          X"0B02043" WHEN IR&CONT = "10000011100" ELSE
          X"0050100" WHEN IR&CONT = "10000100000" ELSE
          X"0004000" WHEN IR&CONT = "10000100001" ELSE
          X"0B01044" WHEN IR&CONT = "10000100010" ELSE
          X"0050100" WHEN IR&CONT = "10000101000" ELSE
          X"0004000" WHEN IR&CONT = "10000101001" ELSE
          X"0B01045" WHEN IR&CONT = "10000101010" ELSE
          X"0050100" WHEN IR&CONT = "10000110000" ELSE
          X"0004000" WHEN IR&CONT = "10000110001" ELSE
          X"0B01046" WHEN IR&CONT = "10000110010" ELSE
          X"0050100" WHEN IR&CONT = "10000111000" ELSE
          X"0004000" WHEN IR&CONT = "10000111001" ELSE
          X"0050100" WHEN IR&CONT = "10000111010" ELSE
          X"0008000" WHEN IR&CONT = "10000111011" ELSE
          X"0B01047" WHEN IR&CONT = "10000111100" ELSE
          X"0050100" WHEN IR&CONT = "10001000000" ELSE
          X"0004000" WHEN IR&CONT = "10001000001" ELSE
          X"0B00848" WHEN IR&CONT = "10001000010" ELSE
          X"0050100" WHEN IR&CONT = "10001001000" ELSE
          X"0004000" WHEN IR&CONT = "10001001001" ELSE
          X"0B00849" WHEN IR&CONT = "10001001010" ELSE
          X"0050100" WHEN IR&CONT = "10001010000" ELSE
          X"0004000" WHEN IR&CONT = "10001010001" ELSE
          X"0B0084A" WHEN IR&CONT = "10001010010" ELSE
          X"0050100" WHEN IR&CONT = "10001011000" ELSE
          X"0004000" WHEN IR&CONT = "10001011001" ELSE
          X"0050100" WHEN IR&CONT = "10001011010" ELSE
          X"0008000" WHEN IR&CONT = "10001011011" ELSE
          X"0B0084B" WHEN IR&CONT = "10001011100" ELSE
          X"0050100" WHEN IR&CONT = "10010000000" ELSE
          X"0004000" WHEN IR&CONT = "10010000001" ELSE
          X"0B82040" WHEN IR&CONT = "10010000010" ELSE
          X"0050100" WHEN IR&CONT = "10010001000" ELSE
          X"0004000" WHEN IR&CONT = "10010001001" ELSE
          X"0B81045" WHEN IR&CONT = "10010001010" ELSE
          X"0050100" WHEN IR&CONT = "10010010000" ELSE
          X"0004000" WHEN IR&CONT = "10010010001" ELSE
          X"0B8084A" WHEN IR&CONT = "10010010010" ELSE
          X"0050100" WHEN IR&CONT = "10010100000" ELSE
          X"0004000" WHEN IR&CONT = "10010100001" ELSE
          X"0C02040" WHEN IR&CONT = "10010100010" ELSE
          X"0050100" WHEN IR&CONT = "10010101000" ELSE
          X"0004000" WHEN IR&CONT = "10010101001" ELSE
          X"0C01045" WHEN IR&CONT = "10010101010" ELSE
          X"0050100" WHEN IR&CONT = "10010110000" ELSE
          X"0004000" WHEN IR&CONT = "10010110001" ELSE
          X"0C0084A" WHEN IR&CONT = "10010110010" ELSE
          X"0050100" WHEN IR&CONT = "10011000000" ELSE
          X"0004000" WHEN IR&CONT = "10011000001" ELSE
          X"0C82040" WHEN IR&CONT = "10011000010" ELSE
          X"0050100" WHEN IR&CONT = "10011001000" ELSE
          X"0004000" WHEN IR&CONT = "10011001001" ELSE
          X"0C81045" WHEN IR&CONT = "10011001010" ELSE
          X"0050100" WHEN IR&CONT = "10011010000" ELSE
          X"0004000" WHEN IR&CONT = "10011010001" ELSE
          X"0C8084A" WHEN IR&CONT = "10011010010" ELSE
          X"0050100" WHEN IR&CONT = "10011111000" ELSE
          X"0804000" WHEN IR&CONT = "10011111001" ELSE
          X"0050100" WHEN IR&CONT = "11001000000" ELSE
          X"0004000" WHEN IR&CONT = "11001000001" ELSE
          X"0D02000" WHEN IR&CONT = "11001000010" ELSE
          X"0050100" WHEN IR&CONT = "11001001000" ELSE
          X"0004000" WHEN IR&CONT = "11001001001" ELSE
          X"0D01004" WHEN IR&CONT = "11001001010" ELSE
          X"0050100" WHEN IR&CONT = "11001010000" ELSE
          X"0004000" WHEN IR&CONT = "11001010001" ELSE
          X"0D00808" WHEN IR&CONT = "11001010010" ELSE
          X"0050100" WHEN IR&CONT = "11001100000" ELSE
          X"0004000" WHEN IR&CONT = "11001100001" ELSE
          X"0D82000" WHEN IR&CONT = "11001100010" ELSE
          X"0050100" WHEN IR&CONT = "11001101000" ELSE
          X"0004000" WHEN IR&CONT = "11001101001" ELSE
          X"0D81004" WHEN IR&CONT = "11001101010" ELSE
          X"0050100" WHEN IR&CONT = "11001110000" ELSE
          X"0004000" WHEN IR&CONT = "11001110001" ELSE
          X"0D80808" WHEN IR&CONT = "11001110010" ELSE
          X"0050100" WHEN IR&CONT = "10100000000" ELSE
          X"0004000" WHEN IR&CONT = "10100000001" ELSE
          X"0900400" WHEN IR&CONT = "10100000010" ELSE
          X"0050100" WHEN IR&CONT = "10100001000" ELSE
          X"0004000" WHEN IR&CONT = "10100001001" ELSE
          X"0900401" WHEN IR&CONT = "10100001010" ELSE
          X"0050100" WHEN IR&CONT = "10100010000" ELSE
          X"0004000" WHEN IR&CONT = "10100010001" ELSE
          X"0900402" WHEN IR&CONT = "10100010010" ELSE
          X"0050100" WHEN IR&CONT = "10100011000" ELSE
          X"0004000" WHEN IR&CONT = "10100011001" ELSE
          X"0050100" WHEN IR&CONT = "10100011010" ELSE
          X"0008000" WHEN IR&CONT = "10100011011" ELSE
          X"0900403" WHEN IR&CONT = "10100011100" ELSE
          X"0050100" WHEN IR&CONT = "10100100000" ELSE
          X"0004000" WHEN IR&CONT = "10100100001" ELSE
          X"0900404" WHEN IR&CONT = "10100100010" ELSE
          X"0050100" WHEN IR&CONT = "10100101000" ELSE
          X"0004000" WHEN IR&CONT = "10100101001" ELSE
          X"0900405" WHEN IR&CONT = "10100101010" ELSE
          X"0050100" WHEN IR&CONT = "10100110000" ELSE
          X"0004000" WHEN IR&CONT = "10100110001" ELSE
          X"0900406" WHEN IR&CONT = "10100110010" ELSE
          X"0050100" WHEN IR&CONT = "10100111000" ELSE
          X"0004000" WHEN IR&CONT = "10100111001" ELSE
          X"0050100" WHEN IR&CONT = "10100111010" ELSE
          X"0008000" WHEN IR&CONT = "10100111011" ELSE
          X"0900407" WHEN IR&CONT = "10100111100" ELSE
          X"0050100" WHEN IR&CONT = "10101000000" ELSE
          X"0004000" WHEN IR&CONT = "10101000001" ELSE
          X"0900408" WHEN IR&CONT = "10101000010" ELSE
          X"0050100" WHEN IR&CONT = "10101001000" ELSE
          X"0004000" WHEN IR&CONT = "10101001001" ELSE
          X"0900409" WHEN IR&CONT = "10101001010" ELSE
          X"0050100" WHEN IR&CONT = "10101010000" ELSE
          X"0004000" WHEN IR&CONT = "10101010001" ELSE
          X"090040A" WHEN IR&CONT = "10101010010" ELSE
          X"0050100" WHEN IR&CONT = "10101011000" ELSE
          X"0004000" WHEN IR&CONT = "10101011001" ELSE
          X"0050100" WHEN IR&CONT = "10101011010" ELSE
          X"0008000" WHEN IR&CONT = "10101011011" ELSE
          X"090040B" WHEN IR&CONT = "10101011100" ELSE
          X"0050100" WHEN IR&CONT = "1011----000" ELSE
          X"0004000" WHEN IR&CONT = "1011----001" ELSE
          X"0050100" WHEN IR&CONT = "1011----010" ELSE
          X"0008000" WHEN IR&CONT = "1011----011" ELSE
          X"0840040" WHEN IR&CONT = "1011----100" ELSE
          X"0050100" WHEN IR&CONT = "11000000000" ELSE
          X"0004000" WHEN IR&CONT = "11000000001" ELSE
          X"0050100" WHEN IR&CONT = "11000000010" ELSE
          X"0008000" WHEN IR&CONT = "11000000011" ELSE
          X"0840000" WHEN IR&CONT = "11000000100" ELSE
          X"0050100" WHEN IR&CONT = "11000001000" ELSE
          X"0004000" WHEN IR&CONT = "11000001001" ELSE
          X"0050100" WHEN IR&CONT = "11000001010" ELSE
          X"0008000" WHEN IR&CONT = "11000001011" ELSE
          X"0840000" WHEN IR&CONT = "11000001100" ELSE
          X"0050100" WHEN IR&CONT = "11000010000" ELSE
          X"0004000" WHEN IR&CONT = "11000010001" ELSE
          X"0050100" WHEN IR&CONT = "11000010010" ELSE
          X"0008000" WHEN IR&CONT = "11000010011" ELSE
          X"0840000" WHEN IR&CONT = "11000010100" ELSE
          X"0050100" WHEN IR&CONT = "11010000000" ELSE
          X"0004000" WHEN IR&CONT = "11010000001" ELSE
          X"0008010" WHEN IR&CONT = "11010000010" ELSE
          X"0010020" WHEN IR&CONT = "11010000011" ELSE
          X"0008000" WHEN IR&CONT = "11010000100" ELSE
          X"0802003" WHEN IR&CONT = "11010000101" ELSE
          X"0050100" WHEN IR&CONT = "11010001000" ELSE
          X"0004000" WHEN IR&CONT = "11010001001" ELSE
          X"0008015" WHEN IR&CONT = "11010001010" ELSE
          X"0010020" WHEN IR&CONT = "11010001011" ELSE
          X"0008000" WHEN IR&CONT = "11010001100" ELSE
          X"0802003" WHEN IR&CONT = "11010001101" ELSE
          X"0050100" WHEN IR&CONT = "11010010000" ELSE
          X"0004000" WHEN IR&CONT = "11010010001" ELSE
          X"000801A" WHEN IR&CONT = "11010010010" ELSE
          X"0010020" WHEN IR&CONT = "11010010011" ELSE
          X"0008000" WHEN IR&CONT = "11010010100" ELSE
          X"0802003" WHEN IR&CONT = "11010010101" ELSE
          X"0050100" WHEN IR&CONT = "11010100000" ELSE
          X"0004000" WHEN IR&CONT = "11010100001" ELSE
          X"0008010" WHEN IR&CONT = "11010100010" ELSE
          X"0010020" WHEN IR&CONT = "11010100011" ELSE
          X"0008000" WHEN IR&CONT = "11010100100" ELSE
          X"0801007" WHEN IR&CONT = "11010100101" ELSE
          X"0050100" WHEN IR&CONT = "11010101000" ELSE
          X"0004000" WHEN IR&CONT = "11010101001" ELSE
          X"0008015" WHEN IR&CONT = "11010101010" ELSE
          X"0010020" WHEN IR&CONT = "11010101011" ELSE
          X"0008000" WHEN IR&CONT = "11010101100" ELSE
          X"0801007" WHEN IR&CONT = "11010101101" ELSE
          X"0050100" WHEN IR&CONT = "11010110000" ELSE
          X"0004000" WHEN IR&CONT = "11010110001" ELSE
          X"000801A" WHEN IR&CONT = "11010110010" ELSE
          X"0010020" WHEN IR&CONT = "11010110011" ELSE
          X"0008000" WHEN IR&CONT = "11010110100" ELSE
          X"0801007" WHEN IR&CONT = "11010110101" ELSE
          X"0050100" WHEN IR&CONT = "11011000000" ELSE
          X"0004000" WHEN IR&CONT = "11011000001" ELSE
          X"0008010" WHEN IR&CONT = "11011000010" ELSE
          X"0010020" WHEN IR&CONT = "11011000011" ELSE
          X"0008000" WHEN IR&CONT = "11011000100" ELSE
          X"080080B" WHEN IR&CONT = "11011000101" ELSE
          X"0050100" WHEN IR&CONT = "11011001000" ELSE
          X"0004000" WHEN IR&CONT = "11011001001" ELSE
          X"0008010" WHEN IR&CONT = "11011001010" ELSE
          X"0010020" WHEN IR&CONT = "11011001011" ELSE
          X"0008000" WHEN IR&CONT = "11011001100" ELSE
          X"080080B" WHEN IR&CONT = "11011001101" ELSE
          X"0050100" WHEN IR&CONT = "11011010000" ELSE
          X"0004000" WHEN IR&CONT = "11011010001" ELSE
          X"0008010" WHEN IR&CONT = "11011010010" ELSE
          X"0010020" WHEN IR&CONT = "11011010011" ELSE
          X"0008000" WHEN IR&CONT = "11011010100" ELSE
          X"080080B" WHEN IR&CONT = "11011010101" ELSE
          X"0050100" WHEN IR&CONT = "11100000000" ELSE
          X"0004000" WHEN IR&CONT = "11100000001" ELSE
          X"0008010" WHEN IR&CONT = "11100000010" ELSE
          X"0010020" WHEN IR&CONT = "11100000011" ELSE
          X"0008010" WHEN IR&CONT = "11100000100" ELSE
          X"0800200" WHEN IR&CONT = "11100000101" ELSE
          X"0050100" WHEN IR&CONT = "11100001000" ELSE
          X"0004000" WHEN IR&CONT = "11100001001" ELSE
          X"0008010" WHEN IR&CONT = "11100001010" ELSE
          X"0010020" WHEN IR&CONT = "11100001011" ELSE
          X"0008015" WHEN IR&CONT = "11100001100" ELSE
          X"0800200" WHEN IR&CONT = "11100001101" ELSE
          X"0050100" WHEN IR&CONT = "11100010000" ELSE
          X"0004000" WHEN IR&CONT = "11100010001" ELSE
          X"0008010" WHEN IR&CONT = "11100010010" ELSE
          X"0010020" WHEN IR&CONT = "11100010011" ELSE
          X"000801A" WHEN IR&CONT = "11100010100" ELSE
          X"0800200" WHEN IR&CONT = "11100010101" ELSE
          X"0050100" WHEN IR&CONT = "11100100000" ELSE
          X"0004000" WHEN IR&CONT = "11100100001" ELSE
          X"0008015" WHEN IR&CONT = "11100100010" ELSE
          X"0010020" WHEN IR&CONT = "11100100011" ELSE
          X"0008010" WHEN IR&CONT = "11100100100" ELSE
          X"0800200" WHEN IR&CONT = "11100100101" ELSE
          X"0050100" WHEN IR&CONT = "11100101000" ELSE
          X"0004000" WHEN IR&CONT = "11100101001" ELSE
          X"0008015" WHEN IR&CONT = "11100101010" ELSE
          X"0010020" WHEN IR&CONT = "11100101011" ELSE
          X"0008015" WHEN IR&CONT = "11100101100" ELSE
          X"0800200" WHEN IR&CONT = "11100101101" ELSE
          X"0050100" WHEN IR&CONT = "11100110000" ELSE
          X"0004000" WHEN IR&CONT = "11100110001" ELSE
          X"0008015" WHEN IR&CONT = "11100110010" ELSE
          X"0010020" WHEN IR&CONT = "11100110011" ELSE
          X"000801A" WHEN IR&CONT = "11100110100" ELSE
          X"0800200" WHEN IR&CONT = "11100110101" ELSE
          X"0050100" WHEN IR&CONT = "11101000000" ELSE
          X"0004000" WHEN IR&CONT = "11101000001" ELSE
          X"000801A" WHEN IR&CONT = "11101000010" ELSE
          X"0010020" WHEN IR&CONT = "11101000011" ELSE
          X"0008010" WHEN IR&CONT = "11101000100" ELSE
          X"0800200" WHEN IR&CONT = "11101000101" ELSE
          X"0050100" WHEN IR&CONT = "11101001000" ELSE
          X"0004000" WHEN IR&CONT = "11101001001" ELSE
          X"000801A" WHEN IR&CONT = "11101001010" ELSE
          X"0010020" WHEN IR&CONT = "11101001011" ELSE
          X"0008015" WHEN IR&CONT = "11101001100" ELSE
          X"0800200" WHEN IR&CONT = "11101001101" ELSE
          X"0050100" WHEN IR&CONT = "11101010000" ELSE
          X"0004000" WHEN IR&CONT = "11101010001" ELSE
          X"000801A" WHEN IR&CONT = "11101010010" ELSE
          X"0010020" WHEN IR&CONT = "11101010011" ELSE
          X"000801A" WHEN IR&CONT = "11101010100" ELSE
          X"0800200" WHEN IR&CONT = "11101010101" ELSE
          X"0050100" WHEN IR&CONT = "1111----000" ELSE
          X"0004000" WHEN IR&CONT = "1111----001" ELSE
          X"0050100" WHEN IR&CONT = "1111----010" ELSE
          X"0008000" WHEN IR&CONT = "1111----011" ELSE
          X"1000000" WHEN IR&CONT = "1111----100" ELSE
          X"0840040" WHEN IR&CONT = "1111----101" ELSE
          X"0050100" WHEN IR&CONT = "10011110000" ELSE
          X"0004000" WHEN IR&CONT = "10011110001" ELSE
          X"0840080" WHEN IR&CONT = "10011110010" ELSE
          X"08700C0";
			 
			 salida_mem_control <= se�ales_de_control(24 downto 0);

end Behavioral;

