library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM is
port (clk : in std_logic;
      rom_enable: in std_logic;
      direccion : in std_logic_vector(9 downto 0);
      rom_datos : out std_logic_vector(7 downto 0));
end ROM;

architecture syn of ROM is
    type rom_type is array (0 to 1023) of std_logic_vector (7 downto 0);                 
    signal ROM : rom_type:= (X"20", X"2C", X"13", X"00", X"20", X"24", X"1C", X"05",
                             X"B0", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                             X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
									  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00");
    
	 signal rdata : std_logic_vector(7 downto 0);
begin

    rdata <= ROM(conv_integer(direccion));

    process (clk)
    begin
        if (clk'event and clk = '1') then
            if (rom_enable = '1') then
                rom_datos <= rdata;
				else
					rom_datos <= "ZZZZZZZZ";
            end if;
        end if;
    end process;

end syn;

				